* AD797 SPICE Macro-model 
* Description: Amplifier
* Generic Desc: 10/30V, BIP, OP, Low THD, Low Noise, 1X
* Developed by: AAG / PMI
* Revision History: 08/10/2012 - Updated to new header style
* 1.0 (10/1992)
* Copyright 1992, 2012 by Analog Devices, Inc.
*
* Refer to http://www.analog.com/Analog_Root/static/techSupport/designTools/spiceModels/license/spice_general.html for License Statement.  Use of this model
* indicates your acceptance with the terms and provisions in the License Statement.
*
* BEGIN Notes:
*
* Not Modeled:
*    
* Parameters modeled include: 
*
* END Notes
*
* Node assignments
*             non-inverting input
*             | inverting input
*             | | positive supply
*             | | |  negative supply
*             | | |  |  output
*             | | |  |  |  decompensation
*             | | |  |  |  |
.SUBCKT AD797 1 2 99 50 38 14
*
* INPUT STAGE & POLE AT 500 MHz
*
IOS 1 2 DC 50E-9
CIND 1 2 20E-12
CINC1 1 98 5E-12
GRCM1 1 98 POLY(2) 1 31 2 31 (0,5E-9,5E-9)
GN1 0 1 44 0 1E-3
CINC2 2 98 5E-12
GRCM2 2 98 POLY(2) 1 31 2 31 (0,5E-9,5E-9)
GN2 0 2 47 0 1E-3
EOS 9 3 POLY(1) 22 31 25E-6 1
EN 3 1 41 0 0.1
D1 2 9 DX
D2 9 2 DX
Q1 5 2 4 QX
Q2 6 9 4 QX
R3 97 5 0.5172
R4 97 6 0.5172
C2 5 6 3.0772E-10
I1 4 51 100E-3
EPOS 97 0 99 0 1
ENEG 51 0 50 0 1
*
* INPUT VOLTAGE NOISE GENERATOR
*
VN1 40 0 DC 2
DN1 40 41 DEN
DN2 41 42 DEN
VN2 0 42 DC 2
*
* +INPUT CURRENT NOISE GENERATOR
*
VN3 43 0 DC 2
DN3 43 44 DIN
DN4 44 45 DIN
VN4 0 45 DC 2
*
* -INPUT CURRENT NOISE GENERATOR
*
VN5 46 0 DC 2
DN5 46 47 DIN
DN6 47 48 DIN
VN6 0 48 DC 2
*
* GAIN STAGE & DOMINANT POLE AT 7.33 Hz
*
EREF 98 0 31 0 1
G1 98 10 5 6 10
R7 10 98 10
E1 99 11 POLY(1) 99 31 -2.294 1
D3 10 11 DX
E2 12 50 POLY(1) 31 50 -2.294 1
D4 12 10 DX
G2 98 13 10 31 1E-3
R8 13 98 10
G3 99 14 98 13 34.558E-3
G4 99 16 98 98 34.558E-3
G5 14 15 15 14 20E-3
G6 16 17 17 14 20E-3
R9 15 18 400
R10 17 18 400
E3 18 98 16 98 1
R11 16 98 4.3406E8
C5 16 98 50E-12
V1 99 19 DC 2.2542
D5 16 19 DX
V2 20 50 DC 2.2542
D6 20 16 DX
RDC 14 98 1E15
*
* COMMON-MODE GAIN NETWORK WITH ZERO AT 1.35 kHz
*
ECM 21 98 POLY(2) 1 31 2 31 (0,158.11E-3,158.11E-3)
RCM1 21 22 1
CCM 21 22 1.1789E-4
RCM2 22 98 1E-6
*
* POLE-ZERO PAIR AT 3.9 MHz/10 MHz
*
GPZ 98 23 16 98 1
RPZ1 23 98 1
RPZ2 23 24 0.63934
CPZ 24 98 24.893E-9
*
* NEGATIVE ZERO AT -300 MHz
*
ENZ 25 98 23 31 1E6
RNZ1 25 26 1
CNZ 25 26 -5.3052E-10
RNZ2 26 98 1E-6
*
* POLE AT 300 MHz
*
GP2 98 27 26 31 1
RP2 27 98 1
CP2 27 98 5.3052E-10
*
* POLE AT 500 MHz
*
GP3 98 28 27 31 1
RP3 28 98 1
CP3 28 98 3.1831E-10
*
* POLE AT 500 MHz
*
GP4 98 29 28 31 1
RP4 29 98 1
CP4 29 98 3.1831E-10
*
* OUTPUT STAGE
*
VW 29 30 DC 0
RDC1 99 31 23.25E3
CDC 31 0 1E-6
RDC2 31 50 23.25E3
GO1 98 32 37 30 25E-3
DO1 32 33 DX
VO1 33 98 DC 0
DO2 34 32 DX
VO2 98 34 DC 0
FDC 99 50 POLY(2) VO1 VO2 7.56E-3 1 1
VSC1 35 37 0.945
DSC1 30 35 DX
VSC2 37 36 0.745
DSC2 36 30 DX
FSC1 37 0 VSC1 1
FSC2 0 37 VSC2 1
GO3 37 99 99 30 25E-3
GO4 50 37 30 50 25E-3
RO1 99 37 40
RO2 37 50 40
LO 37 38 10E-9
*
* MODELS USED
*
.MODEL QX NPN(BF=2E5)
.MODEL DX D(IS=1E-15)
.MODEL DEN D(IS=1E-12 RS=6.3708E3 AF=1 KF=1.59E-15)
.MODEL DIN D(IS=1E-12 RS=474 AF=1 KF=7.816E-15)
.ENDS AD797





